module shift_reg
#(
    parameter SIZE = 8
)
(
    input in, clk,
    output reg out
);
    reg [SIZE-1:0] data;

    always @ (posedge clk)
    begin
        out <= data[SIZE-1];
        data <= {data[SIZE-2:0], in};
    end
endmodule

